module graphics_engine (
    input wire vga_clk,             

    input wire [9:0] pixel_x,       
    input wire [9:0] pixel_y,       
    input wire display_area,        
    input wire [9:0] dino_y,        
    input wire [9:0] obstacle_x1,   
    input wire [9:0] obstacle_x2,   
    input wire game_over,           

    output reg [3:0] red,           
    output reg [3:0] green,         
    output reg [3:0] blue          
);

    localparam OBSTACLE_WIDTH  = 50;
    localparam OBSTACLE_HEIGHT = 150;
    localparam DINO_X          = 50;
    localparam DINO_WIDTH      = 50;
    localparam DINO_HEIGHT     = 100;

    wire pixel_in_obstacle1; 
    wire pixel_in_obstacle2;
    wire in_body; 
    wire in_head; 
    wire in_legs; 
    wire in_tail;
    wire in_eye;
    wire pixel_in_dino;

    // Obstacle boundaries
    assign pixel_in_obstacle1 = (pixel_x >= obstacle_x1) &&
                                (pixel_x <  obstacle_x1 + OBSTACLE_WIDTH) &&
                                (pixel_y >= 480 - OBSTACLE_HEIGHT) &&
                                (pixel_y <  480);

    assign pixel_in_obstacle2 = (pixel_x >= obstacle_x2) &&
                                (pixel_x <  obstacle_x2 + OBSTACLE_WIDTH) &&
                                (pixel_y >= 480 - OBSTACLE_HEIGHT) &&
                                (pixel_y <  480);

    // [generated by CHATGPT because I can't draw]
    assign in_body = (pixel_x >= DINO_X + 10) &&
                     (pixel_x <  DINO_X + 40) &&
                     (pixel_y >= 480 - dino_y - 60) &&
                     (pixel_y <  480 - dino_y);

    assign in_head = (pixel_x >= DINO_X + 35) &&
                     (pixel_x <  DINO_X + 48) &&
                     (pixel_y >= 480 - dino_y - 80) &&
                     (pixel_y <  480 - dino_y - 60);

    assign in_legs = ((pixel_x >= DINO_X + 12 && pixel_x < DINO_X + 18) || 
                      (pixel_x >= DINO_X + 32 && pixel_x < DINO_X + 38)) &&
                     (pixel_y >= 480 - dino_y && pixel_y < 480 - dino_y + 10);

    assign in_tail = (pixel_x >= DINO_X) &&
                     (pixel_x <  DINO_X + 10) &&
                     (pixel_y >= 480 - dino_y - 30) &&
                     (pixel_y <  480 - dino_y + 10);

    assign in_eye  = (pixel_x == DINO_X + 45) &&
                     (pixel_y == 480 - dino_y - 75);

    assign pixel_in_dino = in_body || in_head || in_legs || in_tail || in_eye;

    always @(posedge vga_clk) 
    begin
        if (display_area) 
        begin
            if (pixel_in_obstacle1 || pixel_in_obstacle2 || pixel_in_dino) 
            begin
                red   <= 4'd8;
                green <= 4'd8;
                blue  <= 4'd8;
            end 
            else 
            begin
                red   <= 4'd15;
                green <= 4'd15;
                blue  <= 4'd15;
            end
        end 
        else 
        begin
            red   <= 4'd0;
            green <= 4'd0;
            blue  <= 4'd0;
        end
    end

endmodule
